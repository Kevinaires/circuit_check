library ieee;
use ieee.std_logic_1164.all;

entity NAND_ent is
port(   x: in bit;
        y: in bit;
        F: out bit
);
end NAND_ent;  

--------------------------------------------------

architecture behav1 of NAND_ent is
begin

    process(x, y)
    begin
        -- compare to truth table
        if ((x='1') and (y='1')) then
            F <= '0';
        else
            F <= '1';
        end if;
    end process;

end behav1;