Sorry, no second example yet.
